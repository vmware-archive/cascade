module foo();
endmodule
