module foo#(
  parameter X=10, y=10, z=10, // Comma-separated list of parameters
  parameter W=10)             // Single-element declaration
();
endmodule
