module conds();
  always begin
    if (cond);

    if (cond) begin
    end
  
    if (cond) begin
    end
    else if (cond) begin
    end

    if (cond);
    else begin
    end
  end
endmodule
