module foo(x,y,z);
  input wire x;
  input wire y;
  input wire z;
endmodule
