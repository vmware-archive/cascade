module foo();
  input  wire x1,x2,x3;
  inout  wire y;
  output wire z;
  output reg r1;
  output reg r2,r3=5,r4;
endmodule
