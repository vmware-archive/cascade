module and(x,y,z);
  input wire x;
  input wire y;
  output wire z;

  assign z = x & y;
endmodule
