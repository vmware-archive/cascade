// A module named foo hasn't been declared
foo f();
