reg x[1:0][1:0];
always @(x) begin

end
initial $finish;
