module foo(x, .y(Y));
endmodule
