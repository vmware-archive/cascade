module foo#(
  parameter X=10,Y=20,Z=30 // Single declaration with multiple trailing assignments
)();
endmodule
