module foo();
  initial begin
    w = 10;
    y <= 30;
  end
endmodule
