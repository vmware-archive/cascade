module foo(x);
