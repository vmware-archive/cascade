module foo();
  foo f();
endmodule

initial $finish;
