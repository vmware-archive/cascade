module foo(x, y);
endmodule
