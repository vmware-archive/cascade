module foo();
endmodule

foo f();
initial $finish;
