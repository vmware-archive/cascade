module foo(
    input wire x
  );
  input wire y;
endmodule
