(* w *) (* x, y=1, z="hello" *) module foo();
endmodule
