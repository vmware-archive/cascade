module foo();
  assign x1 = y1;
  assign x2 = y2, x3 = y3;
endmodule
