module foo(
  input wire x,y,z,      // Comma-separated list of inputs
  output wire a,b,c,     // Comma-separated list of outputs
  output reg q=1,s,t=1   // Comma-separated list of outputs with assignments intermixed 
);
endmodule
