genvar i;
always @(posedge clock.val) begin
  if (i) begin end
end
