module foo();
  input wire x;
endmodule
