module foo#(
  parameter X = 10,       
  parameter Y = 20
)(
  input wire x,
  output wire y,
  inout wire z
);

endmodule
