wire x;
always @(posedge clock.val) begin
  x = 1;
end
