module foo();
  initial begin
    $write("Hello ");
    $display("World");
    $finish;
  end
endmodule
