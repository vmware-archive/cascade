// This file has trailing whitespace before the EOF

module foo();
endmodule







